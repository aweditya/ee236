I-V Characteristic of Solar Cell for different levels of illumination

* Include model file
.include ../../../models/lab-4/Solar_Cell.txt

* Netlist
vs 1 0 dc 1 ac 0
r 1 2 100
x 2 0 solar_cell

.control

set temp=35
dc vs -2 2 0.001

meas dc voc find v(2) when i(vs)=0
meas dc isc find i(vs) when v(2)=0
print voc isc

print -i(vs) v(2) > ../results/iv-0-35

set temp=45
dc vs -2 2 0.001

meas dc voc find v(2) when i(vs)=0
meas dc isc find i(vs) when v(2)=0
print voc isc

print -i(vs) v(2) > ../results/iv-0-45

set temp=55
dc vs -2 2 0.001

meas dc voc find v(2) when i(vs)=0
meas dc isc find i(vs) when v(2)=0
print voc isc

print -i(vs) v(2) > ../results/iv-0-55

set temp=65
dc vs -2 2 0.001

meas dc voc find v(2) when i(vs)=0
meas dc isc find i(vs) when v(2)=0
print voc isc

print -i(vs) v(2) > ../results/iv-0-65

set temp=75
dc vs -2 2 0.001

meas dc voc find v(2) when i(vs)=0
meas dc isc find i(vs) when v(2)=0
print voc isc

print -i(vs) v(2) > ../results/iv-0-75

.endc
.end
