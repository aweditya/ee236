Simulation Exercise - IV Characteristic of 1N914

* Include 1N914 model files
.include ../../../../models/diodes/Diode_1N914.txt

* Netlist
vs 1 0 dc 1 ac 0
r1 1 2 100
r2 2 0 1k

v 2 3 dc 0 ac 0
r3 3 4 100
d 4 0 1n914

.dc vs -200 5 0.05
.control
run

plot i(v) vs v(4)
print v(4) i(v) > ../results/1n914

set color0=white
set color1=black
set color2=red
.endc
.end
