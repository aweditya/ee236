Diode I-V Characteristic and Band Gap

* Include LED and Diode model files
.include ../../../models/diodes/Diode_1N914.txt
.include ../../../models/leds/blue_5mm.txt
.include ../../../models/leds/green_5mm.txt
.include ../../../models/leds/red_5mm.txt
.include ../../../models/leds/white_5mm.txt

* Netlist
vs 1 0 dc 1 ac 0

vreg 1 2 dc 0 ac 0
rreg 2 7 100
dreg 7 0 1n914

vblue 1 3 dc 0 ac 0
rblue 3 8 100
dblue 8 0 blue

vgreen 1 4 dc 0 ac 0
rgreen 4 9 100
dgreen 9 0 green 

vred 1 5 dc 0 ac 0
rred 5 10 100
dred 10 0 red

vwhite 1 6 dc 0 ac 0
rwhite 6 11 100
dwhite 11 0 white

.dc vs 0.01 5 0.005
.control
run
meas dc cutoff_regular find v(7) when i(vreg)=1m 
meas dc cutoff_blue find v(8) when i(vblue)=1m 
meas dc cutoff_green find v(9) when i(vgreen)=1m 
meas dc cutoff_red find v(10) when i(vred)=1m 
meas dc cutoff_white find v(11) when i(vwhite)=1m 

plot i(vreg) vs v(7), i(vblue) vs v(8), i(vgreen) vs v(9), i(vred) vs v(10), i(vwhite) vs v(11)
plot ln(i(vreg)) vs v(7), ln(i(vblue)) vs v(8), ln(i(vgreen)) vs v(9), ln(i(vred)) vs v(10), ln(i(vwhite)) vs v(11)

print v(7) i(vreg) > ../results/regularDiode
print v(8) i(vblue) > ../results/blueLED
print v(9) i(vgreen) > ../results/greenLED
print v(10) i(vred) > ../results/redLED
print v(11) i(vwhite) > ../results/whiteLED

.endc
.end
