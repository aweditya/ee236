Bridge Rectifier using BAT85

* Include the diode model file
.include ../../../../models/lab-2/BAT85.txt

* AC source: sin(offset amplitude FREQ delay damping-factor)
vin 1 0 sin(0 5 50 0 0)

* Bridge rectifier
x1 1 2 bat85
x2 3 1 bat85
x3 3 0 bat85
x4 0 2 bat85
rL 2 3 1k

.tran 1us 40ms
.control
run

plot v(1) v(2,3)
plot v(2,3) vs v(1)

set color0=white
set color1=black
set color2=red

print v(1) v(2,3) > ../results/voltage-bat85

.endc
.end
