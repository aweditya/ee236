Simulation Exercise - IV Characteristic of Zener 

* Include zener model files
.include ../../../../models/diodes/Zener_1N4688.txt

* Netlist
vs 1 0 dc 1 ac 0
r1 1 2 100
r2 2 0 1k

v 2 3 dc 0 ac 0
r3 3 4 100
x 4 0 1n4688

.dc vs -200 5 0.05
.control
run

plot i(v) vs v(4)
print v(4) i(v) > ../results/zener

set color0=white
set color1=black
set color2=red
.endc
.end
